library verilog;
use verilog.vl_types.all;
entity sc_interrupt_tb is
end sc_interrupt_tb;
