module flopr(clk, rst, d, q);
  input clk;
  input rst;
  input d;
  output q;
endmodule